`define DATA_IN_WIDTH 8